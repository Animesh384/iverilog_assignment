module bitmutiplexcer(input s0,s1,i0,i1,i2,i3,output f);
    assign f=(~s0&~s1&i0)|(~s0&s1&i1)|(s0&~s1&i2)|(s0&s1&i3);
endmodule