module hello_world;
  initial
  begin
	  $display("hello world");
  end
endmodule
