module test_comparator;
    reg a,b;
    wire g,e,l;
    comparator a1(a,b,g,e,l);
    initial begin
        $dumpfile("gtkwave.vcd");
        $dumpvars;
        $display($time,"time|a|b|g|e|l|");
        $monitor($time,"time|%d|%d|%d|%d|%d|",a,b,g,e,l);
        a=0; b=0;
        #10  a=0; b=1;
        #10  a=1; b=0;
        #10  a=1; b=1;
        #10 $finish;
    end
endmodule